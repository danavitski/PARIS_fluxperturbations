netcdf paris_protocol {
dimensions:
	time = 12 ;
	longitude = 250 ; 
	latitude = 390 ; 
	countrynumber = 43; 
variables:
	int time(time) ;
		time:standard_name = "time" ;
		time:units = "seconds since 2000-01-01T00:00:00Z" ;
		time:calendar = "standard" ;
		time:axis = "T" ;
	double longitude(longitude) ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:axis = "X" ;
	double latitude(latitude) ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:axis = "Y" ;
	float flux_ff_exchange_prior(time, latitude, longitude) ;
		flux_ff_exchange_prior:long_name = "prior anthropogenic CO2 fluxes" ;
		flux_ff_exchange_prior:comment = "" ;
		flux_ff_exchange_prior:dtype = "float" ;
		flux_ff_exchange_prior:units = "mol m-2 s-1" ;
	float flux_ocean_exchange_prior(time, latitude, longitude) ;
		flux_ocean_exchange_prior:long_name = "prior ocean CO2 fluxes" ;
		flux_ocean_exchange_prior:comment = "" ;
		flux_ocean_exchange_prior:dtype = "float" ;
		flux_ocean_exchange_prior:units = "mol m-2 s-1" ;
	float flux_bio_exchange_prior(time, latitude, longitude) ;
		flux_bio_exchange_prior:long_name = "prior biosphere CO2 fluxes" ;
		flux_bio_exchange_prior:comment = "" ;
		flux_bio_exchange_prior:dtype = "float" ;
		flux_bio_exchange_prior:units = "mol m-2 s-1" ;
	float flux_fire_exchange_prior(time, latitude, longitude) ;
		flux_fire_exchange_prior:long_name = "prior wildfire CO2 fluxes" ;
		flux_fire_exchange_prior:comment = "" ;
		flux_fire_exchange_prior:dtype = "float" ;
		flux_fire_exchange_prior:units = "mol m-2 s-1" ;
	float flux_ff_exchange_posterior(time, latitude, longitude) ;
		flux_ff_exchange_posterior:long_name = "posterior anthropogenic CO2 fluxes" ;
		flux_ff_exchange_posterior:comment = "" ;
		flux_ff_exchange_posterior:dtype = "float" ;
		flux_ff_exchange_posterior:units = "mol m-2 s-1" ;
	float flux_ocean_exchange_posterior(time, latitude, longitude) ;
		flux_ocean_exchange_posterior:long_name = "posterior ocean CO2 fluxes" ;
		flux_ocean_exchange_posterior:comment = "" ;
		flux_ocean_exchange_posterior:dtype = "float" ;
		flux_ocean_exchange_posterior:units = "mol m-2 s-1" ;
	float flux_bio_exchange_posterior(time, latitude, longitude) ;
		flux_bio_exchange_posterior:long_name = "posterior biosphere CO2 fluxes" ;
		flux_bio_exchange_posterior:comment = "" ;
		flux_bio_exchange_posterior:dtype = "float" ;
		flux_bio_exchange_posterior:units = "mol m-2 s-1" ;
	float flux_fire_exchange_posterior(time, latitude, longitude) ;
		flux_fire_exchange_posterior:long_name = "posterior wildfire CO2 fluxes" ;
		flux_fire_exchange_posterior:comment = "" ;
		flux_fire_exchange_posterior:dtype = "float" ;
		flux_fire_exchange_posterior:units = "mol m-2 s-1" ;
	float country_flux_ff_posterior(time, countrynumber) ;
		country_flux_ff_exchange_posterior:long_name = "country-averaged posterior fossil fuel CO2 fluxes" ;
		country_flux_ff_exchange_posterior:comment = "" ;
		country_flux_ff_exchange_posterior:dtype = "float" ;
		country_flux_ff_exchange_posterior:units = "mol m-2 s-1" ;
	float country_flux_ocean_exchange_posterior(time, countrynumber) ;
		country_flux_ocean_exchange_posterior:long_name = "country-averaged posterior ocean CO2 fluxes" ;
		country_flux_ocean_exchange_posterior:comment = "" ;
		country_flux_ocean_exchange_posterior:dtype = "float" ;
		country_flux_ocean_exchange_posterior:units = "mol m-2 s-1" ;
	float country_flux_bio_exchange_posterior(time, countrynumber) ;
		country_flux_bio_exchange_posterior:long_name = "country-averaged posterior biosphere CO2 fluxes" ;
		country_flux_bio_exchange_posterior:comment = "" ;
		country_flux_bio_exchange_posterior:dtype = "float" ;
		country_flux_bio_exchange_posterior:units = "mol m-2 s-1" ;
	float country_flux_fire_exchange_posterior(time, countrynumber) ;
		country_flux_fire_exchange_posterior:long_name = "country-averaged posterior wildfire CO2 fluxes" ;
		country_flux_fire_exchange_posterior:comment = "" ;
		country_flux_fire_exchange_posterior:dtype = "float" ;
		country_flux_fire_exchange_posterior:units = "mol m-2 s-1" ;
	float uncertainty_country_flux_ff_prior(time, countrynumber, countrynumber) ;
		uncertainty_country_flux_ff_prior:long_name = "uncertainty matrix of country-averaged prior fossil fuel CO2 fluxes" ;
		uncertainty_country_flux_ff_prior:comment = "" ;
		uncertainty_country_flux_ff_prior:dtype = "float" ;
    	uncertainty_country_flux_ff_prior:units = "mol m-2 s-1" ;
	float uncertainty_country_flux_ocean_prior(time, countrynumber, countrynumber) ;
		uncertainty_country_flux_ocean_prior:long_name = "uncertainty matrix of country-averaged prior ocean CO2 fluxes" ;
		uncertainty_country_flux_ocean_prior:comment = "" ;
		uncertainty_country_flux_ocean_prior:dtype = "float" ;
    	uncertainty_country_flux_ocean_prior:units = "mol m-2 s-1" ;
	float uncertainty_country_flux_bio_prior(time, countrynumber, countrynumber) ;
		uncertainty_country_flux_bio_prior:long_name = "uncertainty matrix of country-averaged prior biosphere CO2 fluxes" ;
		uncertainty_country_flux_bio_prior:comment = "" ;
		uncertainty_country_flux_bio_prior:dtype = "float" ;
    	uncertainty_country_flux_bio_prior:units = "mol m-2 s-1" ;
	float uncertainty_country_flux_fire_prior(time, countrynumber, countrynumber) ;
		uncertainty_country_flux_fire_prior:long_name = "uncertainty matrix of country-averaged prior wildfire CO2 fluxes" ;
		uncertainty_country_flux_fire_prior:comment = "" ;
		uncertainty_country_flux_fire_prior:dtype = "float" ;
    	uncertainty_country_flux_fire_prior:units = "mol m-2 s-1" ;
  	float uncertainty_country_flux_ff_posterior(time, countrynumber, countrynumber) ;
		uncertainty_country_flux_ff_posterior:long_name = "uncertainty matrix of country-averaged posterior fossil fuel CO2 fluxes" ;
		uncertainty_country_flux_ff_posterior:comment = "" ;
		uncertainty_country_flux_ff_posterior:dtype = "float" ;
    	uncertainty_country_flux_ff_posterior:units = "mol m-2 s-1" ;
	float uncertainty_country_flux_ocean_posterior(time, countrynumber, countrynumber) ;
		uncertainty_country_flux_ocean_posterior:long_name = "uncertainty matrix of country-averaged posterior ocean CO2 fluxes" ;
		uncertainty_country_flux_ocean_posterior:comment = "" ;
		uncertainty_country_flux_ocean_posterior:dtype = "float" ;
    	uncertainty_country_flux_ocean_posterior:units = "mol m-2 s-1" ;
	float uncertainty_country_flux_bio_posterior(time, countrynumber, countrynumber) ;
		uncertainty_country_flux_bio_posterior:long_name = "uncertainty matrix of country-averaged posterior biosphere CO2 fluxes" ;
		uncertainty_country_flux_bio_posterior:comment = "" ;
		uncertainty_country_flux_bio_posterior:dtype = "float" ;
    	uncertainty_country_flux_bio_posterior:units = "mol m-2 s-1" ;
	float uncertainty_country_flux_fire_posterior(time, countrynumber, countrynumber) ;
		uncertainty_country_flux_fire_posterior:long_name = "uncertainty matrix of country-averaged posterior wildfire CO2 fluxes" ;
		uncertainty_country_flux_fire_posterior:comment = "" ;
		uncertainty_country_flux_fire_posterior:dtype = "float" ;
    	uncertainty_country_flux_fire_posterior:units = "mol m-2 s-1" ;

// global attributes:
	:summary = "A collection of monthly-averaged CTE-HR CO2 fluxes for 2021, containing hourly estimates of biospheric fluxes, anthropogenic emissions (total and per sector), GFAS fire emissions and Jena CarboScope ocean fluxes, all re-gridded to match the resolution of the biospheric fluxes." ;
	:source = "CTE-HR 1.0. Created using the code from https://git.wageningenur.nl/ctdas/CTDAS/-/tree/near-real-time, hash b8e1a8f" ;
    :model_name = "CarbonTracker Europe - High Resolution" ;
	:frequency = "monthly" ;
	:geospatial_lat_resolution = "0.1 degree" ;
	:geospatial_lon_resolution = "0.2 degree" ;
	:crs = "spherical earth with radius of 6370 km" ;
	:institution = "Wageningen University, department of Meteorology and Air Quality, Wageningen, the Netherlands; \n Rijksuniversiteit Groningen, Groningen, the Netherlands; \n ICOS Carbon Portal, Lund, Sweden" ;
	:contact = "Daan Kivits, Wageningen University & Research, daan.kivits@wur.nl" ;
	:project = "Process Attribution of Regional emISsions (PARIS)"
	:keywords = "carbon flux, carbontracker, emission model, flux product" ;
	:license = "CC-BY-4.0" ;
	:Conventions = "CF-1.8" ;
	:references = "van der Woude et al. (2023), https://doi.org/10.5194/essd-15-579-2023" ;
	:comment = "Positive terrestrial and oceanic biosphere fluxes are emissions, and negative mean uptake. For more information, see https://doi.org/10.5281/zenodo.6477331. The country names that correspond to the given country numbers can be found in the CTE-HR base flux set and accessory country mask file"
	:history = "" ;
}
